<svg viewBox="0 0 250 80" xmlns="http://www.w3.org/2000/svg">
  <!-- خلفية الشعار -->
  <linearGradient id="logoGradient" x1="0%" y1="0%" x2="100%" y2="100%">
    <stop offset="0%" stop-color="#3a7bd5" />
    <stop offset="100%" stop-color="#00d2ff" />
  </linearGradient>
  
  <!-- رمز الأستاذ -->
  <g transform="translate(25, 15)">
    <!-- رمز الكتاب -->
    <path d="M0,0 L40,0 L40,50 L20,40 L0,50 Z" fill="url(#logoGradient)" stroke="#fff" stroke-width="2" />
    <!-- رمز القلم -->
    <path d="M50,10 L55,5 L65,15 L60,20 L50,10 Z M48,12 L20,40 L15,50 L25,45 L53,17 Z" fill="#2c3e50" />
  </g>
  
  <!-- نص الشعار -->
  <g transform="translate(120, 35)">
    <text font-family="'Tajawal', sans-serif" font-size="24" font-weight="700" fill="#2c3e50" text-anchor="middle" alignment-baseline="middle">
      منصة الأساتذة
    </text>
    <text font-family="'Tajawal', sans-serif" font-size="14" font-weight="400" fill="#3a7bd5" text-anchor="middle" alignment-baseline="middle" y="20">
      التعليم بطريقة معاصرة
    </text>
  </g>
</svg>